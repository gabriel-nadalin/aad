module mask(q1, q2, q3, out);
	input [2:0] q1;
   input [2:0] q2;
   input [2:0] q3;
   output [8:0] out;